////////////////////////////////////////////////////////////////////////////////////////////////////

`include "encoder.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps
localparam CLOCK_TICK = 5;
localparam CLOCK_MARGIN = 1;

////////////////////////////////////////////////////////////////////////////////////////////////////

module test();

    logic clk;
    logic rst_n;
    logic [ENC_SYM_NUM - 1 : 0][EGF_ORDER - 1 : 0] data_in;
    logic [2 * ENC_SYM_NUM - 2 : 0][EGF_ORDER - 1 : 0] data_out;
    
    encoder test (
        .clk(clk),
        .rst_n(rst_n),
        .data_in(data_in),
        .data_out(data_out)
    );
    
    initial begin
        clk = 0;
        forever #CLOCK_TICK clk = ~clk;
    end
    
    initial begin
        rst_n <= #(0 * CLOCK_TICK) 0;
        rst_n <= #(21 * CLOCK_TICK + CLOCK_MARGIN) 1;
    end
    
    initial begin
        #(20 * CLOCK_TICK + CLOCK_MARGIN);
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(2 * CLOCK_TICK) data_in = '{4'b0000, 4'b0001, 4'b0010, 4'b0011};
        #(2 * CLOCK_TICK) data_in = '{4'b0100, 4'b0101, 4'b0110, 4'b0111};
        #(2 * CLOCK_TICK) data_in = '{4'b1000, 4'b1001, 4'b1010, 4'b1011};
        #(2 * CLOCK_TICK) data_in = '{4'b1100, 4'b1101, 4'b1110, 4'b1111};
        #(100 * CLOCK_TICK) $finish;
    end

//    initial begin
//        #(20 * CLOCK_TICK + CLOCK_MARGIN);
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(2 * CLOCK_TICK) data_in = '{5'b00000, 5'b00001, 5'b00010, 5'b00011, 5'b00100, 5'b00101, 5'b00110, 5'b00111};
//        #(2 * CLOCK_TICK) data_in = '{5'b01000, 5'b01001, 5'b01010, 5'b01011, 5'b01100, 5'b01101, 5'b01110, 5'b01111};
//        #(2 * CLOCK_TICK) data_in = '{5'b10000, 5'b10001, 5'b10010, 5'b10011, 5'b10100, 5'b10101, 5'b10110, 5'b10111};
//        #(2 * CLOCK_TICK) data_in = '{5'b11000, 5'b11001, 5'b11010, 5'b11011, 5'b11100, 5'b11101, 5'b11110, 5'b11111};
//        #(100 * CLOCK_TICK) $finish;
//    end

endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////