////////////////////////////////////////////////////////////////////////////////////////////////////

`include "encoder.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////

module enc_controller (
    input clk,
    input rst_n,
    output logic [$clog2(RS_COD_LEN) - 1 : 0] con_master_counter
);

////////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk) begin
        if (!rst_n) begin
            con_master_counter <= '0;
        end else if (con_master_counter + ENC_SYM_NUM > RS_COD_LEN) begin
            con_master_counter <= con_master_counter + ENC_SYM_NUM - RS_COD_LEN;
        end else begin
            con_master_counter <= con_master_counter + ENC_SYM_NUM;
        end
    end

endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////